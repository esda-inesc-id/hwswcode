// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXIL_MACC_TESTER_MWRAP_MEM_NO_READ_ON_WRITE 0
// Core Configuration Macros.
`define IOB_AXIL_MACC_TESTER_MWRAP_ADDR_W 32
`define IOB_AXIL_MACC_TESTER_MWRAP_DATA_W 32
`define IOB_AXIL_MACC_TESTER_MWRAP_INIT_MEM 1
`define IOB_AXIL_MACC_TESTER_MWRAP_USE_INTMEM 1
`define IOB_AXIL_MACC_TESTER_MWRAP_MEM_ADDR_W 18
`define IOB_AXIL_MACC_TESTER_MWRAP_FW_BASEADDR 0
`define IOB_AXIL_MACC_TESTER_MWRAP_FW_ADDR_W 18
`define IOB_AXIL_MACC_TESTER_MWRAP_RST_POL 1
`define IOB_AXIL_MACC_TESTER_MWRAP_BOOTROM_ADDR_W 12
// Core Constants. DO NOT CHANGE
`define IOB_AXIL_MACC_TESTER_MWRAP_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_AXIL_MACC_TESTER_MWRAP_AXI_ID_W 1
`define IOB_AXIL_MACC_TESTER_MWRAP_AXI_ADDR_W 18
`define IOB_AXIL_MACC_TESTER_MWRAP_AXI_DATA_W 32
`define IOB_AXIL_MACC_TESTER_MWRAP_AXI_LEN_W 4
`define IOB_AXIL_MACC_TESTER_MWRAP_BOOTROM_MEM_HEXFILE "iob_axil_macc_tester_bootrom"
`define IOB_AXIL_MACC_TESTER_MWRAP_EXT_MEM_HEXFILE "iob_axil_macc_tester_firmware"
