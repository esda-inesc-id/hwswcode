// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXIL_MACC_CSRS_DATA_W 32
// Core Constants. DO NOT CHANGE
`define IOB_AXIL_MACC_CSRS_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_AXIL_MACC_CSRS_ADDR_W 4
