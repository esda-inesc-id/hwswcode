// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define IOB_TIMER_CORE_VERSION 16'h0081
