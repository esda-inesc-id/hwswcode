// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXIL_MACC_TESTER_IOB_VEXRISCV_AXI_ID_W 0
`define IOB_AXIL_MACC_TESTER_IOB_VEXRISCV_AXI_ADDR_W 0
`define IOB_AXIL_MACC_TESTER_IOB_VEXRISCV_AXI_DATA_W 0
`define IOB_AXIL_MACC_TESTER_IOB_VEXRISCV_AXI_LEN_W 0
// Core Constants. DO NOT CHANGE
`define IOB_AXIL_MACC_TESTER_IOB_VEXRISCV_VERSION 16'h0001
