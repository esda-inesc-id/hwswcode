// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXIL_MACC_TESTER_AXI_FULL_XBAR_MERGE_ID_W 1
`define IOB_AXIL_MACC_TESTER_AXI_FULL_XBAR_MERGE_LEN_W 1
// Core Constants. DO NOT CHANGE
`define IOB_AXIL_MACC_TESTER_AXI_FULL_XBAR_MERGE_VERSION 16'h0081
