`timescale 1ns / 1ps
`include "iob_axil_macc_tester_syn_conf.vh"

module iob_axil_macc_tester_syn (
);


endmodule
