// general_operation: General operation group
// Core Configuration Macros.
`define IOB_AXIL_MACC_TESTER_ADDR_W 32
`define IOB_AXIL_MACC_TESTER_DATA_W 32
`define IOB_AXIL_MACC_TESTER_INIT_MEM 1
`define IOB_AXIL_MACC_TESTER_USE_INTMEM 1
`define IOB_AXIL_MACC_TESTER_MEM_ADDR_W 18
`define IOB_AXIL_MACC_TESTER_FW_BASEADDR 0
`define IOB_AXIL_MACC_TESTER_FW_ADDR_W 18
`define IOB_AXIL_MACC_TESTER_RST_POL 1
`define IOB_AXIL_MACC_TESTER_BOOTROM_ADDR_W 12
// Core Constants. DO NOT CHANGE
`define IOB_AXIL_MACC_TESTER_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_AXIL_MACC_TESTER_AXI_ID_W 1
`define IOB_AXIL_MACC_TESTER_AXI_ADDR_W 18
`define IOB_AXIL_MACC_TESTER_AXI_DATA_W 32
`define IOB_AXIL_MACC_TESTER_AXI_LEN_W 4
`define IOB_AXIL_MACC_TESTER_BOOTROM_MEM_HEXFILE "iob_axil_macc_tester_bootrom"
`define IOB_AXIL_MACC_TESTER_EXT_MEM_HEXFILE "iob_axil_macc_tester_firmware"
