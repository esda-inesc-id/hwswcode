// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define IOB_AXIL2IOB_VERSION 16'h0081
