// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_TIMER_CSRS_DATA_W 32
`define IOB_TIMER_CSRS_WDATA_W 1
// Core Constants. DO NOT CHANGE
`define IOB_TIMER_CSRS_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_TIMER_CSRS_ADDR_W 4
